
// Module: ModuleKeyword
module ModuleKeyword ();
endmodule

// Module: MacroModuleKeyword
macromodule MacroModuleKeyword ();
endmodule

// Module: StaticLifetime
module static StaticLifetime ();
endmodule

// Module: AutomaticLifetime
module automatic AutomaticLifetime ();
endmodule

// Module: Complex_Identifier$
module Complex_Identifier$ ();
endmodule

// Module: NamedEnd
module NamedEnd ();
endmodule: NamedEnd

// Module: NamedEnd_Complex_Identifier$
module NamedEnd_Complex_Identifier$ ();
endmodule: NamedEnd_Complex_Identifier$
