
// Group: 1-1 Modules
//

// Module: Module11A
module Module11A #(int x) (int y);
endmodule

// Module: Module11B
module Module11B #(int xx) (int y);
endmodule

// Module: Module11C
module Module11C #(int x) (int yy);
endmodule

// Module: Module11D
module Module11D #(int x) ();
endmodule

// Module: Module11E
module Module11E #() (int y);
endmodule


// Group: 2-1 Modules
//

// Module: Module21A
module Module21A #(int x, int y) (int z);
endmodule

// Module: Module21B
module Module21B #(int xx, int y) (int z);
endmodule

// Module: Module21C
module Module21C #(int x, int yy) (int z);
endmodule

// Module: Module21D
module Module21D #(int x, int y) (int zz);
endmodule

// Module: Module21E
module Module21E #(int x, int y) ();
endmodule

// Module: Module21F
module Module21F #(int xx, int y) ();
endmodule

// Module: Module21G
module Module21G #(int x, int yy) ();
endmodule


// Group: 1-2 Modules
//

// Module: Module12A
module Module12A #(int x) (int y, int z);
endmodule

// Module: Module12B
module Module12B #(int xx) (int y, int z);
endmodule

// Module: Module12C
module Module12C #(int x) (int yy, int z);
endmodule

// Module: Module12D
module Module12D #(int x) (int y, int zz);
endmodule

// Module: Module12E
module Module12E #() (int y, int z);
endmodule

// Module: Module12F
module Module12F #() (int yy, int z);
endmodule

// Module: Module12G
module Module12G #() (int y, int zz);
endmodule
