
/*
	Topic: Strings

		--- code ---

		simple = "abc def";

		embeddedQuotes = "int \" int \" int";

		backslashTrap1 = "abc\\";

		backslashTrap2 = "int \\\" int \\\" int";

		escapedLineBreak = "abc \
		def";

		---

*/