
/*
	Topic: Keywords

		--- code ---

		module  // keyword

		always_latch  // keyword with underscore

		supply1  // keyword with number

		Module  // identifier, keywords must be lowercase

		MODULE  // identifier, keywords must be lowercase

		_module  // identifier

		$module  // identifier

		\module  // escaped identifer, not a keyword

		\(module)  // escaped identifiers continue until whitespace, not a keyword

		some_module  // identifier

		some$module  // identifiers can have $ characters

		module$  // identifier

		module_  // identifier

		$error  // keyword

		error // identifier

		$error_  // identifier

		$$error  // identifier

		x$error  // identifier

		_$error  // identifier

		---
*/